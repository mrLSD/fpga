`define NUMBER_1 'b11000000 
`define NUMBER_2 'b11000000
`ifndef NUMBER_3
	`define NUMBER_3 'b11000000
`endif 