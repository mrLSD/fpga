`define NUMBER_0 'b11000000 
`define NUMBER_1 'b11111001
`define NUMBER_2 'b10100100
`define NUMBER_3 'b10110000
`define NUMBER_4 'b10011001
`define NUMBER_5 'b10010010
`define NUMBER_6 'b10000010
`define NUMBER_7 'b11111000
`define NUMBER_8 'b10000000
`define NUMBER_9 'b10010000

`define DIGIT_BLOCK_1 6'b111110
`define DIGIT_BLOCK_2 6'b111101
`define DIGIT_BLOCK_3 6'b111011
`define DIGIT_BLOCK_4 6'b110111
`define DIGIT_BLOCK_5 6'b101111
`define DIGIT_BLOCK_6 6'b011111
`define DIGIT_BLOCK_EMPTY 6'b111111

`define DIGIT_COUNT_LIMIT 30000
//`define CLOCK_TIME_LIMIT 26'h2_FFF_F00
`define CLOCK_TIME_LIMIT 50_000_000
