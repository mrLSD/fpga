package fonts;

parameter reg [0:7] FONT1 [0:1] [0:63] = '{
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf8, 8'h3f, 8'hfc, 8'h70, 8'h0e, 8'h67, 8'he6, 8'h6f, 8'hf6, 8'h6c, 8'h36, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h36, 8'h6f, 8'hf6, 8'h67, 8'he6, 8'h70, 8'h0e, 8'h3f, 8'hfc, 8'h1f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 0 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}   /* 1 */
};
//module get_font_16x32();
endpackage