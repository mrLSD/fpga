module vga(
   clock,
   switch,
   disp_RGB,
   hsync,
   vsync
);
parameter string tst = "SystemVerilog";
wire [0:15] arr1 [0:255] [0:63] = '{
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf8, 8'h3f, 8'hfc, 8'h70, 8'h0e, 8'h67, 8'he6, 8'h6f, 8'hf6, 8'h6c, 8'h36, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h06, 8'h6c, 8'h36, 8'h6f, 8'hf6, 8'h67, 8'he6, 8'h70, 8'h0e, 8'h3f, 8'hfc, 8'h1f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 0 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 1 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 2 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h07, 8'he0, 8'h07, 8'he0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 3 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h03, 8'hc0, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h3f, 8'hfc, 8'h7f, 8'hfe, 8'h7f, 8'hfe, 8'h3f, 8'hfc, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 4 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf8, 8'h3f, 8'hf8, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 5 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'hf8, 8'h0f, 8'hf8, 8'h1c, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3f, 8'hfc, 8'h7f, 8'hfe, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00},  /* 6 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hc0, 8'h07, 8'he0, 8'h07, 8'he0, 8'h07, 8'he0, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 7 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1d, 8'hb8, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h1d, 8'hb8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 8 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h07, 8'hf8, 8'h07, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 9 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h30, 8'h3c, 8'h30, 8'h7c, 8'h30, 8'hec, 8'h31, 8'hcc, 8'h33, 8'h8c, 8'h37, 8'h0c, 8'h3e, 8'h0c, 8'h3c, 8'h0c, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 10 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h30, 8'h3c, 8'h30, 8'h7c, 8'h30, 8'hec, 8'h31, 8'hcc, 8'h33, 8'h8c, 8'h37, 8'h0c, 8'h3e, 8'h0c, 8'h3c, 8'h0c, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 11 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hfc, 8'h07, 8'hfc, 8'h0e, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h1c, 8'h0c, 8'h38, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 12 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 13 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h1f, 8'hf8, 8'h1f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 14 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0e, 8'h1f, 8'hff, 8'h0f, 8'hff, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h00},  /* 15 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 16 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h8c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 17 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h8c, 8'h1f, 8'hfe, 8'h0f, 8'hff, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h00},  /* 18 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hf0, 8'h00, 8'hf0, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h38, 8'h3f, 8'hf0, 8'h3f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 19 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hfc, 8'h3f, 8'hfc, 8'h71, 8'h8c, 8'h61, 8'h8c, 8'h61, 8'h8c, 8'h61, 8'h8c, 8'h61, 8'h8c, 8'h61, 8'h8c, 8'h71, 8'h8c, 8'h3f, 8'h8c, 8'h1f, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 20 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h1c, 8'h38, 8'h18, 8'h18, 8'h18, 8'h00, 8'h1c, 8'h00, 8'h0f, 8'hc0, 8'h0f, 8'he0, 8'h18, 8'h70, 8'h18, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h1c, 8'h18, 8'h0e, 8'h18, 8'h07, 8'hf0, 8'h03, 8'hf0, 8'h00, 8'h38, 8'h00, 8'h18, 8'h18, 8'h18, 8'h1c, 8'h38, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 21 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h7f, 8'h0c, 8'h7f, 8'h8c, 8'h61, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h61, 8'hcc, 8'h7f, 8'h8c, 8'h7f, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 22 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h38, 8'h3f, 8'hf0, 8'h3f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 23 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h03, 8'hc0, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h1d, 8'hb8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 24 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1d, 8'hb8, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 25 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h70, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h7f, 8'hfe, 8'h7f, 8'hfe, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h00, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 26 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h7f, 8'hfe, 8'h7f, 8'hfe, 8'h38, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 27 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h07, 8'hfc, 8'h07, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 28 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'hf0, 8'h61, 8'hf8, 8'h63, 8'h9c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h7f, 8'h0c, 8'h7f, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h9c, 8'h61, 8'hf8, 8'h60, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 29 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'hec, 8'h01, 8'hcc, 8'h03, 8'h8c, 8'h07, 8'h0c, 8'h0e, 8'h0c, 8'h1c, 8'h0c, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 30 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf0, 8'h38, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 31 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 32 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 33 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 34 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 35 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h80, 8'h31, 8'h80, 8'h31, 8'h80, 8'h39, 8'h80, 8'h1f, 8'hf0, 8'h0f, 8'hf8, 8'h01, 8'h9c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 36 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1e, 8'h18, 8'h3f, 8'h18, 8'h33, 8'h30, 8'h33, 8'h30, 8'h3f, 8'h60, 8'h1e, 8'h60, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h00, 8'h03, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h0c, 8'hf0, 8'h0d, 8'hf8, 8'h19, 8'h98, 8'h19, 8'h98, 8'h31, 8'hf8, 8'h30, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 37 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'h80, 8'h1f, 8'hc0, 8'h38, 8'he0, 8'h30, 8'h60, 8'h30, 8'h60, 8'h30, 8'h60, 8'h38, 8'he0, 8'h1d, 8'hc0, 8'h0f, 8'h80, 8'h0f, 8'h00, 8'h1f, 8'h8c, 8'h39, 8'hdc, 8'h70, 8'hf8, 8'h60, 8'h70, 8'h60, 8'h30, 8'h60, 8'h30, 8'h60, 8'h70, 8'h70, 8'hf8, 8'h3f, 8'hdc, 8'h1f, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 38 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 39 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h03, 8'h00, 8'h07, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h07, 8'h00, 8'h03, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 40 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'he0, 8'h00, 8'hc0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 41 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h38, 8'h38, 8'h1c, 8'h70, 8'h0e, 8'he0, 8'h07, 8'hc0, 8'h03, 8'h80, 8'h7f, 8'hfc, 8'h7f, 8'hfc, 8'h03, 8'h80, 8'h07, 8'hc0, 8'h0e, 8'he0, 8'h1c, 8'h70, 8'h38, 8'h38, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 42 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 43 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h80, 8'h03, 8'h00, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 44 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 45 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 46 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h00, 8'h03, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 47 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h30, 8'h3c, 8'h30, 8'h7c, 8'h30, 8'hec, 8'h31, 8'hcc, 8'h33, 8'h8c, 8'h37, 8'h0c, 8'h3e, 8'h0c, 8'h3c, 8'h0c, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 48 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h03, 8'h80, 8'h07, 8'h80, 8'h0f, 8'h80, 8'h0d, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h0f, 8'hf0, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 49 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 50 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h07, 8'hf8, 8'h07, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 51 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h00, 8'h3c, 8'h00, 8'h7c, 8'h00, 8'hec, 8'h01, 8'hcc, 8'h03, 8'h8c, 8'h07, 8'h0c, 8'h0e, 8'h0c, 8'h1c, 8'h0c, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 52 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 53 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf8, 8'h1f, 8'hf8, 8'h38, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 54 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h00, 8'h18, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 55 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 56 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h1f, 8'hf8, 8'h1f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 57 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 58 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h80, 8'h03, 8'h00, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 59 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h70, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 60 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 61 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h70, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 62 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 63 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf0, 8'h3f, 8'hf8, 8'h70, 8'h1c, 8'h60, 8'h0c, 8'h61, 8'hfc, 8'h63, 8'hfc, 8'h67, 8'h0c, 8'h66, 8'h0c, 8'h66, 8'h0c, 8'h66, 8'h0c, 8'h66, 8'h0c, 8'h66, 8'h0c, 8'h66, 8'h0c, 8'h67, 8'h1c, 8'h63, 8'hfc, 8'h61, 8'hec, 8'h60, 8'h00, 8'h70, 8'h00, 8'h3f, 8'hfc, 8'h1f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 64 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 65 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h3f, 8'hf0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 66 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 67 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hc0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h18, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h30, 8'h38, 8'h3f, 8'hf0, 8'h3f, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 68 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 69 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 70 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'hfc, 8'h30, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 71 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 72 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'he0, 8'h07, 8'he0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 73 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7e, 8'h00, 8'h7e, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h38, 8'h38, 8'h1f, 8'hf0, 8'h0f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 74 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h30, 8'h38, 8'h30, 8'h70, 8'h30, 8'he0, 8'h31, 8'hc0, 8'h33, 8'h80, 8'h37, 8'h00, 8'h3e, 8'h00, 8'h3c, 8'h00, 8'h3c, 8'h00, 8'h3e, 8'h00, 8'h37, 8'h00, 8'h33, 8'h80, 8'h31, 8'hc0, 8'h30, 8'he0, 8'h30, 8'h70, 8'h30, 8'h38, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 75 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 76 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h70, 8'h1c, 8'h78, 8'h3c, 8'h6c, 8'h6c, 8'h6c, 8'h6c, 8'h67, 8'hcc, 8'h63, 8'h8c, 8'h63, 8'h8c, 8'h61, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 77 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h3c, 8'h0c, 8'h3e, 8'h0c, 8'h37, 8'h0c, 8'h33, 8'h8c, 8'h31, 8'hcc, 8'h30, 8'hec, 8'h30, 8'h7c, 8'h30, 8'h3c, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 78 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 79 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 80 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h31, 8'hcc, 8'h38, 8'hfc, 8'h1f, 8'hf8, 8'h0f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 81 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h37, 8'h00, 8'h33, 8'h80, 8'h31, 8'hc0, 8'h30, 8'he0, 8'h30, 8'h70, 8'h30, 8'h38, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 82 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h00, 8'h1f, 8'hf0, 8'h0f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 83 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 84 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 85 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 86 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h61, 8'h0c, 8'h63, 8'h8c, 8'h63, 8'h8c, 8'h67, 8'hcc, 8'h6c, 8'h6c, 8'h6c, 8'h6c, 8'h78, 8'h3c, 8'h70, 8'h1c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 87 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h06, 8'h60, 8'h06, 8'h60, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h06, 8'h60, 8'h06, 8'h60, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h18, 8'h18, 8'h18, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 88 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h06, 8'h60, 8'h06, 8'h60, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 89 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 90 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'he0, 8'h0f, 8'he0, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0f, 8'he0, 8'h0f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 91 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 92 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'he0, 8'h0f, 8'he0, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'h0f, 8'he0, 8'h0f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 93 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h03, 8'hc0, 8'h07, 8'he0, 8'h0e, 8'h70, 8'h1c, 8'h38, 8'h38, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 94 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 95 */
    '{8'h00, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 96 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf0, 8'h1f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 97 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 98 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 99 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 100 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 101 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7e, 8'h00, 8'hfe, 8'h01, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h1f, 8'hf8, 8'h1f, 8'hf8, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 102 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h1f, 8'hf8, 8'h1f, 8'hf0, 8'h00, 8'h00},  /* 103 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 104 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h80, 8'h07, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 105 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h78, 8'h00, 8'h78, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h1c, 8'h38, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h00, 8'h00},  /* 106 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h1c, 8'h18, 8'h38, 8'h18, 8'h70, 8'h18, 8'he0, 8'h19, 8'hc0, 8'h1b, 8'h80, 8'h1f, 8'h00, 8'h1f, 8'h00, 8'h1b, 8'h80, 8'h19, 8'hc0, 8'h18, 8'he0, 8'h18, 8'h70, 8'h18, 8'h38, 8'h18, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 107 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h80, 8'h07, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 108 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h31, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 109 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 110 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 111 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf8, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00},  /* 112 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h00},  /* 113 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h33, 8'hfc, 8'h37, 8'hfc, 8'h3e, 8'h00, 8'h3c, 8'h00, 8'h38, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 114 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h00, 8'h1f, 8'hf0, 8'h0f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 115 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h3f, 8'hf0, 8'h3f, 8'hf0, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h80, 8'h01, 8'hfc, 8'h00, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 116 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 117 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 118 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 119 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1c, 8'h38, 8'h0e, 8'h70, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h03, 8'hc0, 8'h07, 8'he0, 8'h0e, 8'h70, 8'h1c, 8'h38, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 120 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h1f, 8'hf8, 8'h1f, 8'hf0, 8'h00, 8'h00},  /* 121 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 122 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hf0, 8'h01, 8'hf0, 8'h03, 8'h80, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h1e, 8'h00, 8'h1e, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h80, 8'h01, 8'hf0, 8'h00, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 123 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 124 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1e, 8'h00, 8'h1f, 8'h00, 8'h03, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'hf0, 8'h00, 8'hf0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h80, 8'h1f, 8'h00, 8'h1e, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 125 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0e, 8'h0c, 8'h1f, 8'h0c, 8'h3b, 8'h8c, 8'h31, 8'hdc, 8'h30, 8'hf8, 8'h30, 8'h70, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 126 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hc0, 8'h3f, 8'he0, 8'h30, 8'h70, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h70, 8'h3f, 8'he0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h3f, 8'hf8, 8'h3f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 127 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 128 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 129 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 130 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h1f, 8'hf8, 8'h1f, 8'hf0, 8'h00, 8'h00},  /* 131 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf0, 8'h1f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 132 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1d, 8'hb8, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h1d, 8'hb8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 133 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h1c, 8'h03, 8'hf8, 8'h03, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 134 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 135 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h07, 8'he0, 8'h03, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 136 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 137 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h1c, 8'h18, 8'h38, 8'h18, 8'h70, 8'h18, 8'he0, 8'h19, 8'hc0, 8'h1b, 8'h80, 8'h1f, 8'h00, 8'h1f, 8'h00, 8'h1b, 8'h80, 8'h19, 8'hc0, 8'h18, 8'he0, 8'h18, 8'h70, 8'h18, 8'h38, 8'h18, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 138 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h80, 8'h07, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 139 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hfc, 8'h07, 8'hfc, 8'h0e, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h1c, 8'h0c, 8'h38, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 140 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h0c, 8'h70, 8'h1c, 8'h78, 8'h3c, 8'h7c, 8'h7c, 8'h6e, 8'hec, 8'h67, 8'hcc, 8'h63, 8'h8c, 8'h61, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 141 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 142 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 143 */
    '{8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 144 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 145 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 146 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 147 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 148 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfe, 8'h0f, 8'hff, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h00},  /* 149 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 150 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h8c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 151 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h8c, 8'h1f, 8'hfe, 8'h0f, 8'hff, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h03, 8'h00, 8'h00},  /* 152 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 153 */
    '{8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 154 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3c, 8'h00, 8'h3c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0f, 8'hf0, 8'h0f, 8'hf8, 8'h0c, 8'h1c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h1c, 8'h0f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 155 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'he0, 8'h07, 8'hf0, 8'h0e, 8'h38, 8'h0c, 8'h18, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h3f, 8'he0, 8'h3f, 8'he0, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h0c, 8'h0c, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 156 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h60, 8'h0c, 8'h7f, 8'h0c, 8'h7f, 8'h8c, 8'h61, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h60, 8'hcc, 8'h61, 8'hcc, 8'h7f, 8'h8c, 8'h7f, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 157 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h1f, 8'he0, 8'h1f, 8'hf0, 8'h18, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h38, 8'h1f, 8'hf0, 8'h1f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 158 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h03, 8'hfc, 8'h03, 8'hfc, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 159 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf0, 8'h1f, 8'hf8, 8'h00, 8'h1c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 160 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h80, 8'h07, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 161 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'hf0, 8'h61, 8'hf8, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h7f, 8'h0c, 8'h7f, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h63, 8'h0c, 8'h61, 8'hf8, 8'h60, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 162 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hfc, 8'h1f, 8'hfc, 8'h38, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h1f, 8'hfc, 8'h0f, 8'hfc, 8'h00, 8'hec, 8'h01, 8'hcc, 8'h03, 8'h8c, 8'h07, 8'h0c, 8'h0e, 8'h0c, 8'h1c, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 163 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h30, 8'h00, 8'h3f, 8'hc0, 8'h3f, 8'hc0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 164 */
    '{8'h00, 8'h00, 8'h0f, 8'h18, 8'h1b, 8'h98, 8'h19, 8'hd8, 8'h18, 8'hf0, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h3c, 8'h0c, 8'h3e, 8'h0c, 8'h37, 8'h0c, 8'h33, 8'h8c, 8'h31, 8'hcc, 8'h30, 8'hec, 8'h30, 8'h7c, 8'h30, 8'h3c, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 165 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 166 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 167 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hf0, 8'h07, 8'hf8, 8'h0e, 8'h1c, 8'h1c, 8'h0e, 8'h38, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'hff, 8'hc0, 8'hff, 8'hc0, 8'h30, 8'h00, 8'h30, 8'h00, 8'hff, 8'hc0, 8'hff, 8'hc0, 8'h30, 8'h00, 8'h30, 8'h00, 8'h38, 8'h00, 8'h1c, 8'h0e, 8'h0e, 8'h1c, 8'h07, 8'hf8, 8'h03, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 168 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc0, 8'h00, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 169 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 170 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h18, 8'h06, 8'h18, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 171 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h60, 8'h18, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 172 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h18, 8'h60, 8'h18, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 173 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'hce, 8'h03, 8'h9c, 8'h07, 8'h38, 8'h0e, 8'h70, 8'h1c, 8'he0, 8'h39, 8'hc0, 8'h73, 8'h80, 8'h73, 8'h80, 8'h39, 8'hc0, 8'h1c, 8'he0, 8'h0e, 8'h70, 8'h07, 8'h38, 8'h03, 8'h9c, 8'h01, 8'hce, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 174 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h73, 8'h80, 8'h39, 8'hc0, 8'h1c, 8'he0, 8'h0e, 8'h70, 8'h07, 8'h38, 8'h03, 8'h9c, 8'h01, 8'hce, 8'h01, 8'hce, 8'h03, 8'h9c, 8'h07, 8'h38, 8'h0e, 8'h70, 8'h1c, 8'he0, 8'h39, 8'hc0, 8'h73, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 175 */
    '{8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00, 8'haa, 8'haa, 8'h00, 8'h00},  /* 176 */
    '{8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55, 8'haa, 8'haa, 8'h55, 8'h55},  /* 177 */
    '{8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa, 8'hff, 8'hff, 8'haa, 8'haa},  /* 178 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 179 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 180 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 181 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hfe, 8'h60, 8'hfe, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 182 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'he0, 8'hff, 8'he0, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 183 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 184 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hfe, 8'h60, 8'hfe, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'hfe, 8'h60, 8'hfe, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 185 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 186 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'he0, 8'hff, 8'he0, 8'h00, 8'h60, 8'h00, 8'h60, 8'hfe, 8'h60, 8'hfe, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 187 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hfe, 8'h60, 8'hfe, 8'h60, 8'h00, 8'h60, 8'h00, 8'h60, 8'hff, 8'he0, 8'hff, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 188 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hff, 8'he0, 8'hff, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 189 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 190 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'h80, 8'hff, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 191 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 192 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 193 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 194 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 195 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 196 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'hff, 8'hff, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 197 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 198 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h7f, 8'h06, 8'h7f, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 199 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h7f, 8'h06, 8'h7f, 8'h06, 8'h00, 8'h06, 8'h00, 8'h07, 8'hff, 8'h07, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 200 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'hff, 8'h07, 8'hff, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h7f, 8'h06, 8'h7f, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 201 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hfe, 8'h7f, 8'hfe, 8'h7f, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 202 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'hfe, 8'h7f, 8'hfe, 8'h7f, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 203 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h7f, 8'h06, 8'h7f, 8'h06, 8'h00, 8'h06, 8'h00, 8'h06, 8'h7f, 8'h06, 8'h7f, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 204 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 205 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hfe, 8'h7f, 8'hfe, 8'h7f, 8'h00, 8'h00, 8'h00, 8'h00, 8'hfe, 8'h7f, 8'hfe, 8'h7f, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 206 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 207 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 208 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 209 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 210 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h07, 8'hff, 8'h07, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 211 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 212 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 213 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'hff, 8'h07, 8'hff, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 214 */
    '{8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'hff, 8'hff, 8'hff, 8'hff, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60, 8'h06, 8'h60},  /* 215 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'hff, 8'hff, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'hff, 8'hff, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 216 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'hff, 8'h80, 8'hff, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 217 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'hff, 8'h01, 8'hff, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 218 */
    '{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff},  /* 219 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff},  /* 220 */
    '{8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00},  /* 221 */
    '{8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff, 8'h00, 8'hff},  /* 222 */
    '{8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 223 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf8, 8'h3f, 8'hfc, 8'h70, 8'h0e, 8'h6f, 8'he6, 8'h6f, 8'hf6, 8'h6c, 8'h36, 8'h6c, 8'h36, 8'h6c, 8'h36, 8'h6f, 8'he6, 8'h6f, 8'hc6, 8'h6d, 8'hc6, 8'h6c, 8'he6, 8'h6c, 8'h76, 8'h70, 8'h0e, 8'h3f, 8'hfc, 8'h1f, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 224 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'he0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h30, 8'h3f, 8'hf0, 8'h3f, 8'hf0, 8'h30, 8'h38, 8'h30, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h0c, 8'h3c, 8'h1c, 8'h37, 8'hf8, 8'h33, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 225 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 226 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 227 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7e, 8'h82, 8'h7e, 8'hc6, 8'h18, 8'hfe, 8'h18, 8'hd6, 8'h18, 8'hc6, 8'h18, 8'hc6, 8'h18, 8'hc6, 8'h18, 8'hc6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 228 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1c, 8'h00, 8'h38, 8'h7f, 8'hfc, 8'h7f, 8'hfc, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h7f, 8'hfc, 8'h7f, 8'hfc, 8'h38, 8'h00, 8'h70, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 229 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h1c, 8'h30, 8'h3c, 8'h30, 8'h7c, 8'h3f, 8'hec, 8'h3f, 8'hcc, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00},  /* 230 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h1f, 8'hf8, 8'h1f, 8'hf8, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 231 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h39, 8'h9c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h39, 8'h9c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 232 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h1f, 8'hf8, 8'h1f, 8'hf8, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h1f, 8'hf8, 8'h1f, 8'hf8, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 233 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc1, 8'h80, 8'hc1, 8'h9c, 8'hc1, 8'hbe, 8'he1, 8'hb6, 8'he1, 8'hb6, 8'hf1, 8'hbe, 8'hf1, 8'h9c, 8'hf9, 8'h80, 8'hd9, 8'h80, 8'hdd, 8'h80, 8'hcd, 8'h80, 8'hcf, 8'h80, 8'hc7, 8'h80, 8'hc7, 8'hbe, 8'hc3, 8'hbe, 8'hc3, 8'h80, 8'hc1, 8'hbe, 8'hc1, 8'hbe, 8'hc1, 8'h80, 8'hc1, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 234 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h31, 8'h8c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 235 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7f, 8'hfc, 8'h7f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 236 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h70, 8'h1c, 8'h38, 8'h38, 8'h1c, 8'h70, 8'h0e, 8'he0, 8'h07, 8'hc0, 8'h03, 8'h80, 8'h03, 8'h80, 8'h07, 8'hc0, 8'h0e, 8'he0, 8'h1c, 8'h70, 8'h38, 8'h38, 8'h70, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 237 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1c, 8'h30, 8'h3e, 8'h30, 8'h36, 8'h60, 8'h36, 8'h60, 8'h3e, 8'hc0, 8'h1c, 8'hc0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h03, 8'h00, 8'h03, 8'h00, 8'h06, 8'h00, 8'h06, 8'h00, 8'h0c, 8'h00, 8'h0c, 8'h00, 8'h19, 8'hdc, 8'h1b, 8'hfe, 8'h33, 8'h76, 8'h33, 8'h76, 8'h63, 8'hfe, 8'h61, 8'hdc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 238 */
    '{8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 239 */
    '{8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h07, 8'he0, 8'h07, 8'he0, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h07, 8'he0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 240 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 241 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h70, 8'h00, 8'h38, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 242 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h38, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0e, 8'h00, 8'h1c, 8'h00, 8'h1c, 8'h00, 8'h0e, 8'h00, 8'h07, 8'h00, 8'h03, 8'h80, 8'h01, 8'hc0, 8'h00, 8'he0, 8'h00, 8'h70, 8'h00, 8'h38, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 243 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hf8, 8'h01, 8'hfc, 8'h01, 8'h8c, 8'h01, 8'h8c, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80},  /* 244 */
    '{8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h31, 8'h80, 8'h31, 8'h80, 8'h3f, 8'h80, 8'h1f, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 245 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3f, 8'hfc, 8'h3f, 8'hfc, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 246 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'h0c, 8'h3f, 8'h9c, 8'h39, 8'hfc, 8'h30, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'h0c, 8'h3f, 8'h9c, 8'h39, 8'hfc, 8'h30, 8'hf8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 247 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'he0, 8'h0f, 8'hf0, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0f, 8'hf0, 8'h07, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 248 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h80, 8'h07, 8'hc0, 8'h07, 8'hc0, 8'h07, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 249 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h01, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 250 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1e, 8'h00, 8'h1e, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h00, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h30, 8'h18, 8'h38, 8'h18, 8'h1c, 8'h18, 8'h0e, 8'h18, 8'h07, 8'h18, 8'h03, 8'h98, 8'h01, 8'hd8, 8'h00, 8'hf8, 8'h00, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 251 */
    '{8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h0f, 8'hf0, 8'h1f, 8'hf8, 8'h38, 8'h1c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 252 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'hc0, 8'h0f, 8'he0, 8'h0c, 8'h60, 8'h0c, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h07, 8'h00, 8'h0f, 8'he0, 8'h0f, 8'he0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 253 */
    '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h1f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00},  /* 254 */
    '{8'h00, 8'h00, 8'h00, 8'h70, 8'h00, 8'he0, 8'h01, 8'hc0, 8'h03, 8'h80, 8'h00, 8'h00, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h30, 8'h0c, 8'h38, 8'h1c, 8'h1f, 8'hf8, 8'h0f, 8'hf0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00}   /* 255 */
};

input  clock;     
input  [1:0]switch;
output [2:0]disp_RGB;
output  hsync;     
output  vsync;     

reg [9:0] hcount;
reg [9:0] vcount;
reg [2:0] data;
reg [2:0] h_dat;
reg [2:0] v_dat;

wire [9:0] x_coord;
wire [9:0] y_coord;

wire  hcount_ov;
wire  vcount_ov;
wire  dat_act;
wire  hsync;
wire  vsync;
reg   vga_clk;

parameter hsync_end   = 10'd95,
   hdat_begin  = 10'd143,
   hdat_end  = 10'd783,
   hpixel_end  = 10'd799,
   vsync_end  = 10'd1,
   vdat_begin  = 10'd34,
   vdat_end  = 10'd514,
   vline_end  = 10'd524;


always @(posedge clock)
begin
 vga_clk = ~vga_clk;
end

always @(posedge vga_clk)
begin
 if (hcount_ov)
  hcount <= 10'd0;
 else
  hcount <= hcount + 10'd1;
end
assign hcount_ov = (hcount == hpixel_end);

always @(posedge vga_clk)
begin
 if (hcount_ov)
 begin
  if (vcount_ov)
   vcount <= 10'd0;
  else
   vcount <= vcount + 10'd1;
 end
end
assign  vcount_ov = (vcount == vline_end);

assign dat_act =    ((hcount >= hdat_begin) && (hcount < hdat_end))
     && ((vcount >= vdat_begin) && (vcount < vdat_end));
assign hsync = (hcount > hsync_end);
assign vsync = (vcount > vsync_end);
assign disp_RGB = (dat_act) ?  data : 3'h00;       

assign x_coord = (hcount - hdat_begin + 1);
assign y_coord = (vcount - vdat_begin + 1);

always @(posedge vga_clk)
begin
 case(switch[1:0])
  2'd0: data <= h_dat;
  2'd1: data <= v_dat;
  2'd2: data <= (v_dat ^ h_dat);
  2'd3: data <= h_dat;
//  2'd3: data <= (v_dat ~^ h_dat);
 endcase
end

always @(posedge vga_clk)
begin
 if((x_coord >= 60 && x_coord < 140) &&
 	(y_coord >= 40 && y_coord < 60) ||
 	(x_coord >= 60 && x_coord < 80) &&
 	(y_coord >= 40 && y_coord < 200) ||
 	(x_coord >= 120 && x_coord < 140) &&
 	(y_coord >= 40 && y_coord < 200) ||
 	(x_coord >= 60 && x_coord < 140) &&
 	(y_coord >= 180 && y_coord < 200)
 	) 
	v_dat <= 3'h6;   
 else 
	v_dat <= 3'h0;
end

wire [9:0]charXPosition;
wire [9:0]charYPosition;
wire [9:0]bitXPosition;
wire [9:0]bitYPosition;

assign charXPosition = (x_coord / 16);
assign charYPosition = (y_coord / 32); 
assign bitXPosition = (x_coord % 16);
assign bitYPosition = (y_coord % 32);

always @(posedge vga_clk)
begin
	h_dat <= 3'h0;
	
	if (charXPosition == 2 && 
		charYPosition == 3
	) begin
		if (arr1[0][bitYPosition][bitXPosition]) begin
			h_dat <= 3'h3;
		end
	end
end

endmodule
