module debouncer(
	input clk, button,
	output reg key_press
);
	
endmodule
